// STAGE 2: INSTRUCTION DECODE UNIT:
// Will generate the Data signals to be delivered to ALU
// Houses the register which may be modified in the write back stage
// Control signals in this unit include RegWrite
 
module Instruction_Decode(clk, reset, Instruction_Code, RegWrite, Write_Data, Write_Register_Num, Read_Data_1, Read_Data_2, Gen_Imm_Data);

//Declaration of inputs of the decode unit
input clk;
input reset;
input [7:0]Instruction_Code; // from the Instruction Fetch Unit; will be connected later
input RegWrite; //will be generated by the control unit
input [7:0] Write_Data; //will be generated during the write back stage
input [2:0] Write_Register_Num;

// Declaration of outputs of the decode unit
output [7:0] Read_Data_1;
output [7:0] Read_Data_2;
output [7:0]Gen_Imm_Data;

// internal connections in the instruction decode segment
wire [2:0]Read_Register_1;
wire [2:0]Read_Register_2;
wire [2:0]Write_Register;

//Assign appropriate bits as per the rs1, rs2 and rd fields to the intermediary wires
assign Read_Register_1=Instruction_Code[5:3];
assign Read_Register_2=Instruction_Code[2:0];

//Generate immediate Data
assign Gen_Imm_Data[7:0] = Instruction_Code[2:0];

// Instantiate the Register file
Register_file RF(Read_Register_1, Read_Register_2, Write_Register_Num, Write_Data, RegWrite, clk, reset, Read_Data_1, Read_Data_2);

endmodule